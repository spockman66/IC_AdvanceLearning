module iic_slave (

    //global clock
    clk,
    rst_n,
    
    iic_scl,
    iic_sda



);


// ----------------port------------------ 
input clk               ;
input rst_n             ;
inout iic_scl           ;
inout iic_sda           ;


// ----------------reg------------------ 
reg []          ;



// ----------------wire------------------ 




// ----------------always------------------ 






// ------------ state machine ----------------- 







endmodule